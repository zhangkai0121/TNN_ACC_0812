`define Tm                              8
`define Tn                              4
`define FEATURE_WIDTH                   24
`define BIAS_WIDTH                      24
`define SCALER_WIDTH                    24
`define KERNEL_WIDTH                    2
`define KERNEL_SIZE                     5
`define FEATURE_SIZE                    28